

module Data_Path_Top_tb;

// Signal Declaration 
    // Common Inputs 
    reg clock;
    reg reset;

// Control Signals
    reg Local_reset;
    
    reg Wr_En_x, Wr_En_A, Wr_En_B, Wr_En_C, Wr_En_D, Wr_En_X;  
    reg Rd_En_x, Rd_En_A, Rd_En_B, Rd_En_C, Rd_En_D, Rd_En_X;
    reg [2:0] MAC_IN_Sel;

    reg [2:0] ROMW_add;
    
    reg [2:0] Sel_Mapping;
    
    // Data Flow
    reg [2*16*16-1:0] Data_In;
    
    wire [2*16*16-1:0] Data_Out;
    
    // Status Signals
    wire Overflow;
    
    integer counter;
    
    // Instantiation
    Data_Path_Top DPUT( 
    .clock(clock),
    .reset(reset),
    .Local_reset(Local_reset),
    .Wr_En_x(Wr_En_x), .Wr_En_A(Wr_En_A), .Wr_En_B(Wr_En_B),
    .Wr_En_C(Wr_En_C), .Wr_En_D(Wr_En_D), .Wr_En_X(Wr_En_X),  
    .Rd_En_x(Rd_En_x), .Rd_En_A(Rd_En_A), .Rd_En_B(Rd_En_B),
    .Rd_En_C(Rd_En_C), .Rd_En_D(Rd_En_D), .Rd_En_X(Rd_En_X),
    .MAC_IN_Sel(MAC_IN_Sel),
    .ROMW_add(ROMW_add),
    .Sel_Mapping(Sel_Mapping),
    .Data_In(Data_In),
    .Data_Out(Data_Out),
    .Overflow(Overflow) 
    );
    
       initial
        begin
        $dumpfile("Data_Path.vcd");
        $dumpvars;
        #1500  $stop ;
        end 
        ///////////initialize inputs 
        initial
        begin
            clock=0;
            reset=0;
            counter=0;
        end
        ///Clock Generator - 100MHZ (10ns Timeperiod)
        initial 
        begin
            clock = 1'b0;
            forever #5 clock= ~clock ;
        end 
        //apply RST to block
        initial
        begin 
        reset = 1'b0;
        #1
        reset = 1'b1;
        #1
        reset = 1'b0;
        #1 ;
        end
        ///////////////////////
        always @(posedge clock)
        begin     
        if(counter == 0)
        begin // reset state
            Local_reset=1;
            Wr_En_x=0;
            Wr_En_A=0;
            Wr_En_B=0;
            Wr_En_C=0; 
            Wr_En_D=0; 
            Wr_En_X=0;  
            Rd_En_x=0;
            Rd_En_A=0; 
            Rd_En_B=0; 
            Rd_En_C=0; 
            Rd_En_D=0; 
            Rd_En_X=0;
            MAC_IN_Sel=3'b000;
            ROMW_add=3'b000;
            Sel_Mapping=3'b000;
            Data_In=512'b00000111_10000001_00001100_00010000_00000100_00000101_00000111_00000001_10000011_10000010_00010000_10000111_00000100_10001001_00000100_10001110_10001111_00000001_10000100_00000010_10000011_00000110_00000001_00001100_00000110_00000100_10001011_10000001_10001111_10000011_00001000_00000011_10001010_10000010_00000010_00001000_00001001_00001011_10000100_00001101_10001000_00000101_00000010_10000100_00001001_10000100_00000010_10000010_00000001_10000100_00001001_00000001_10010000_10000101_00001010_10001000_00001000_10000001_00000011_10000100_10000110_00000101_00000001_10001000 ; 
            counter = counter + 1;
        end
        
         else if(counter == 1)
         begin // Load_x state
            Local_reset = 1'b0;
            Wr_En_x = 1'b1;
            Wr_En_A = 1'b0; 
            Wr_En_B = 1'b0; 
            Wr_En_C = 1'b0;
            Wr_En_D = 1'b0; 
            Wr_En_X = 1'b0; 
            Rd_En_x = 1'b0; 
            Rd_En_A = 1'b0;
            Rd_En_B = 1'b0;
            Rd_En_C = 1'b0;
            Rd_En_D = 1'b0;
            Rd_En_X = 1'b0;
            MAC_IN_Sel  = 3'b000;
            ROMW_add    = 3'b000;       
            Sel_Mapping = 3'b000;
            Data_In= 512'b00000111_10000001_00001100_00010000_00000100_00000101_00000111_00000001_10000011_10000010_00010000_10000111_00000100_10001001_00000100_10001110_10001111_00000001_10000100_00000010_10000011_00000110_00000001_00001100_00000110_00000100_10001011_10000001_10001111_10000011_00001000_00000011_10001010_10000010_00000010_00001000_00001001_00001011_10000100_00001101_10001000_00000101_00000010_10000100_00001001_10000100_00000010_10000010_00000001_10000100_00001001_00000001_10010000_10000101_00001010_10001000_00001000_10000001_00000011_10000100_10000110_00000101_00000001_10001000 ; 
            counter = counter+1;
         end
         else if (counter == 2)
           begin // Load_A State
            Local_reset = 1'b0;
            Wr_En_x = 1'b0;
            Wr_En_A = 1'b1; 
            Wr_En_B = 1'b0; 
            Wr_En_C = 1'b0;
            Wr_En_D = 1'b0; 
            Wr_En_X = 1'b0; 
            Rd_En_x = 1'b1; 
            Rd_En_A = 1'b0;
            Rd_En_B = 1'b0;
            Rd_En_C = 1'b0;
            Rd_En_D = 1'b0;
            Rd_En_X = 1'b0;
            MAC_IN_Sel  = 3'b001;
            ROMW_add    = 3'b001;       
            Sel_Mapping = 3'b001;
            Data_In= 512'b00000111_10000001_00001100_00010000_00000100_00000101_00000111_00000001_10000011_10000010_00010000_10000111_00000100_10001001_00000100_10001110_10001111_00000001_10000100_00000010_10000011_00000110_00000001_00001100_00000110_00000100_10001011_10000001_10001111_10000011_00001000_00000011_10001010_10000010_00000010_00001000_00001001_00001011_10000100_00001101_10001000_00000101_00000010_10000100_00001001_10000100_00000010_10000010_00000001_10000100_00001001_00000001_10010000_10000101_00001010_10001000_00001000_10000001_00000011_10000100_10000110_00000101_00000001_10001000 ; 
            counter = counter+1;
           end
         else if(counter == 3)
         begin //Load_B state
            Local_reset = 1'b0;
            Wr_En_x = 1'b0;
            Wr_En_A = 1'b0; 
            Wr_En_B = 1'b1; 
            Wr_En_C = 1'b0;
            Wr_En_D = 1'b0; 
            Wr_En_X = 1'b0; 
            Rd_En_x = 1'b0; 
            Rd_En_A = 1'b1;
            Rd_En_B = 1'b0;
            Rd_En_C = 1'b0;
            Rd_En_D = 1'b0;
            Rd_En_X = 1'b0;
            MAC_IN_Sel  = 3'b010;
            ROMW_add    = 3'b010;       
            Sel_Mapping = 3'b010;
            Data_In= 512'b00000111_10000001_00001100_00010000_00000100_00000101_00000111_00000001_10000011_10000010_00010000_10000111_00000100_10001001_00000100_10001110_10001111_00000001_10000100_00000010_10000011_00000110_00000001_00001100_00000110_00000100_10001011_10000001_10001111_10000011_00001000_00000011_10001010_10000010_00000010_00001000_00001001_00001011_10000100_00001101_10001000_00000101_00000010_10000100_00001001_10000100_00000010_10000010_00000001_10000100_00001001_00000001_10010000_10000101_00001010_10001000_00001000_10000001_00000011_10000100_10000110_00000101_00000001_10001000 ; 
            counter = counter+1;
         end
         
         else if(counter == 4)
         begin // Load_C state
            Local_reset = 1'b0;
            Wr_En_x = 1'b0;
            Wr_En_A = 1'b0; 
            Wr_En_B = 1'b0; 
            Wr_En_C = 1'b1;
            Wr_En_D = 1'b0; 
            Wr_En_X = 1'b0; 
            Rd_En_x = 1'b0; 
            Rd_En_A = 1'b0;
            Rd_En_B = 1'b1;
            Rd_En_C = 1'b0;
            Rd_En_D = 1'b0;
            Rd_En_X = 1'b0;
            MAC_IN_Sel  = 3'b011;
            ROMW_add    = 3'b011;       
            Sel_Mapping = 3'b011;
            Data_In= 512'b00000111_10000001_00001100_00010000_00000100_00000101_00000111_00000001_10000011_10000010_00010000_10000111_00000100_10001001_00000100_10001110_10001111_00000001_10000100_00000010_10000011_00000110_00000001_00001100_00000110_00000100_10001011_10000001_10001111_10000011_00001000_00000011_10001010_10000010_00000010_00001000_00001001_00001011_10000100_00001101_10001000_00000101_00000010_10000100_00001001_10000100_00000010_10000010_00000001_10000100_00001001_00000001_10010000_10000101_00001010_10001000_00001000_10000001_00000011_10000100_10000110_00000101_00000001_10001000 ; 
            counter = counter+1;
         end
         else if(counter == 5)
         begin // Load_D state
            Local_reset = 1'b0;
            Wr_En_x = 1'b0;
            Wr_En_A = 1'b0; 
            Wr_En_B = 1'b0; 
            Wr_En_C = 1'b0;
            Wr_En_D = 1'b1; 
            Wr_En_X = 1'b0; 
            Rd_En_x = 1'b0; 
            Rd_En_A = 1'b0;
            Rd_En_B = 1'b0;
            Rd_En_C = 1'b1;
            Rd_En_D = 1'b0;
            Rd_En_X = 1'b0;
            MAC_IN_Sel  = 3'b100;
            ROMW_add    = 3'b100;       
            Sel_Mapping = 3'b100;
            Data_In=512'b00000111_10000001_00001100_00010000_00000100_00000101_00000111_00000001_10000011_10000010_00010000_10000111_00000100_10001001_00000100_10001110_10001111_00000001_10000100_00000010_10000011_00000110_00000001_00001100_00000110_00000100_10001011_10000001_10001111_10000011_00001000_00000011_10001010_10000010_00000010_00001000_00001001_00001011_10000100_00001101_10001000_00000101_00000010_10000100_00001001_10000100_00000010_10000010_00000001_10000100_00001001_00000001_10010000_10000101_00001010_10001000_00001000_10000001_00000011_10000100_10000110_00000101_00000001_10001000 ; 
            counter = counter+1;
         end
         
         else if(counter == 6)
         begin // Load_X state
            Local_reset = 1'b0;
            Wr_En_x = 1'b0;
            Wr_En_A = 1'b0; 
            Wr_En_B = 1'b0; 
            Wr_En_C = 1'b0;
            Wr_En_D = 1'b0; 
            Wr_En_X = 1'b1; 
            Rd_En_x = 1'b0; 
            Rd_En_A = 1'b0;
            Rd_En_B = 1'b0;
            Rd_En_C = 1'b0;
            Rd_En_D = 1'b1;
            Rd_En_X = 1'b0;
            MAC_IN_Sel  = 3'b101;
            ROMW_add    = 3'b101;       
            Sel_Mapping = 3'b101;
            Data_In= 512'b00000111_10000001_00001100_00010000_00000100_00000101_00000111_00000001_10000011_10000010_00010000_10000111_00000100_10001001_00000100_10001110_10001111_00000001_10000100_00000010_10000011_00000110_00000001_00001100_00000110_00000100_10001011_10000001_10001111_10000011_00001000_00000011_10001010_10000010_00000010_00001000_00001001_00001011_10000100_00001101_10001000_00000101_00000010_10000100_00001001_10000100_00000010_10000010_00000001_10000100_00001001_00000001_10010000_10000101_00001010_10001000_00001000_10000001_00000011_10000100_10000110_00000101_00000001_10001000 ; 
            counter = counter+1;
         end
         
        end
endmodule    